// `default_nettype none
//
// module buffer(
//     input wire i_clk,
//     input wire i_w_en,
//     input wire[19:0] i_w_data,
//     input wire o_r_en,
//     output wire[19:0] o_w_data
// );
//     reg [3:0] read_addr;
//     reg [3:0] write_addr;
//     reg [19:0] memory [10];
// endmodule
